----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:07:34 10/25/2018 
-- Design Name: 
-- Module Name:    ext - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ext is
    Port ( imm : in  STD_LOGIC_VECTOR (15 downto 0);
           EOp : in  STD_LOGIC_VECTOR (1 downto 0);
           ext : out  STD_LOGIC_VECTOR (31 downto 0));
end ext;

architecture Behavioral of ext is

begin


end Behavioral;

