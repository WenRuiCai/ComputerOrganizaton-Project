`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:25:07 09/25/2018 
// Design Name: 
// Module Name:    MD 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MD(
    input clk,
    input reset,
    input [15:0] D1,
    input [15:0] D2,
    input Start,
    input [0:0] Busy,
    output [15:0] HI,
    output [15:0] LO,
    input MD
    );


endmodule
