`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    22:51:29 11/26/2018
// Design Name:
// Module Name:    Level_WriteBack
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module Level_WriteBack(
    input [31:0] Instr_in,
	 input judge,
    input [31:0] pc_add_4_in,
    input [31:0] pc_add_8_in,
    input [31:0] ALUResult,
    input [31:0] DM_data_in,
    input [4:0] WriteRegNum,
    output [4:0] GRF_A3,
    output WE3,
    output [31:0] Write_GRF_Data
    );

    reg [4:0] Mem_to_Reg=0;
    reg store_WE3=0;

    assign GRF_A3 = WriteRegNum;
    assign WE3 = store_WE3;

    assign Write_GRF_Data=(WriteRegNum==0)?0:((Mem_to_Reg==0)?ALUResult:(
                          (Mem_to_Reg==1)?DM_data_in:pc_add_8_in));

    always @(*) begin
        case (Instr_in[31:26])      //special
            6'b001101:      //ori
                begin
                    Mem_to_Reg=0;
                    store_WE3=1;
                end
            6'b001111:      //lui
                begin
                    Mem_to_Reg=0;
                    store_WE3=1;
                end
            6'b000100:      // beq
                begin
                    Mem_to_Reg=0;
                    store_WE3=0;
                end
				6'b011000:      // blezals
                begin
                    Mem_to_Reg=2;
                    store_WE3=(judge==1)?1:0;
                end
            6'b100011:      //lw
                begin
                    Mem_to_Reg=1;
                    store_WE3=1;
                end
            6'b101011:      //sw
                begin
                    Mem_to_Reg=0;
                    store_WE3=0;
                end
            6'b000011:      //jal
                begin
                    Mem_to_Reg=2;
                    store_WE3=1;
                end
				6'b000010:      //j
                begin
                    Mem_to_Reg=2;
                    store_WE3=0;
                end
            6'b000000:
                begin
                    case (Instr_in[5:0])
                        6'b100001:      //addu
                            begin
                               Mem_to_Reg=0;
                               store_WE3=1;
                            end
                        6'b100011:      //subu
                            begin
                                Mem_to_Reg=0;
                                store_WE3=1;
                            end
                        6'b001000:      //jr
                            begin
                                Mem_to_Reg=0;
                                store_WE3=0;
                            end
                        6'b000000:      //nop
                            begin
                                Mem_to_Reg=0;
                                store_WE3=0;
                            end
                    endcase
                end
        endcase
    end

endmodule
