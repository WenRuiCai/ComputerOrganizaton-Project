`timescale 1ns / 1ps
`include "ALU.v"
`include "mult_and_div.v"
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    22:48:29 11/26/2018
// Design Name:
// Module Name:    Level_Execute
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module Level_Execute(
    input IRQ_E,
    input [6:2] ExcCode_D,
	 input clk,
	 input reset,
    input [31:0] Instr_in,
    input [31:0] PC_plus_4,
    input [31:0] PC_plus_8,
    input [4:0] A1,
    input [4:0] A2,
    input [4:0] A3,
    input [31:0] ReadData1,
    input [31:0] ReadData2,
    input [31:0] ext,
    input [31:0] Data_out_W,
    input [31:0] ALUResult_M,
    input [31:0] jal_pc_from_M,
    input [4:0] select_rs_or_SrcA,
    input [4:0] select_rt_or_SrcB,
    input [31:0] data_from_cp0,
    output [4:0] WriteRegNum,
    output [31:0] rt_value,
    output [31:0] ALUResult_and_HILO,
    output start_mult_div,
	 output busy,
     output WE_cp0,
     output [6:2] ExcCode_E
    );

    wire [31:0] SrcA,SrcB;
    wire [31:0] ALUResult;
    wire [4:0] ALUOp;
    wire [2:0] ALUSrc;

	 wire [31:0] HI,LO;

    reg [4:0] Reg_ALUOP=0;
    reg [2:0] Reg_ALUSrc=0;

    reg [4:0] RegDst=0;

    assign ALUOp = Reg_ALUOP;
	 assign ALUSrc = Reg_ALUSrc;

    assign SrcA=(A1==0)?0:((select_rs_or_SrcA==0)?ReadData1:(
                (select_rs_or_SrcA==1)?ALUResult_M:(
                (select_rs_or_SrcA==2)?Data_out_W:jal_pc_from_M)));

    assign rt_value=(A2==0)?0:((select_rt_or_SrcB==0)?ReadData2:(
                (select_rt_or_SrcB==1)?ALUResult_M:(
                (select_rt_or_SrcB==2)?Data_out_W:jal_pc_from_M)));

    assign SrcB=(ALUSrc==0)?rt_value:ext;

    assign ALUResult_and_HILO = ({Instr_in[31:26]}==6'b000000&&(({Instr_in[5:0]}==6'b010000)))?HI:
                                (({Instr_in[31:26]}==6'b000000&&(({Instr_in[5:0]}==6'b010010)))?LO:
                                (({Instr_in[31:26]}==6'b010000&&{Instr_in[25:21]==5'b00000})?data_from_cp0:ALUResult));

    assign WriteRegNum=(RegDst==0)?A2:(
                       (RegDst==1)?A3:31);

    assign WE_cp0 = ({Instr_in[31:26]}==6'b010000&&{Instr_in[25:21]==5'b00100})?1:0;

    ALU ALU (SrcA,SrcB,Instr_in[10:6],ALUOp,ALUResult);

	 mult_and_div mult_and_div	(clk,reset,IRQ_E,Instr_in,SrcA,rt_value,HI,LO,start_mult_div,busy);

//**************************judge overflow*******************************************//
    integer i=0;
    reg [32:0] judgenumber=0;
    assign ExcCode_E = (i==0)?ExcCode_D:12;
    always @(*) begin
        if({Instr_in[31:26]}==6'b001000||({Instr_in[31:26]}==6'b000000&&{Instr_in[5:0]}==6'b100000)) begin         //add or addi
            judgenumber=$signed(SrcA)+$signed(SrcB);
            if(($signed(judgenumber)>0&&$signed(ALUResult)<=0)||($signed(judgenumber)<0&&$signed(ALUResult)>=0))
                i=1;
            else
                i=0;
        end
        else if({Instr_in[31:26]}==6'b000000&&{Instr_in[5:0]}==6'b100010) begin
            judgenumber=$signed(SrcA)-$signed(SrcB);
            if(($signed(judgenumber)>0&&$signed(ALUResult)<=0)||($signed(judgenumber)<0&&$signed(ALUResult)>=0))
                i=1;
            else
                i=0;
        end
        else
            i=0;
    end
//**************************judge overflow*******************************************//

    /////////////////////////////////////////////////ALUOP ??ALUSrc???
    always @(*) begin
        case (Instr_in[31:26])    //Special
        6'b001101:      //ori
            begin
                Reg_ALUOP=1;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b001110:      //xori
            begin
                Reg_ALUOP=3;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b001100:      //andi
            begin
                Reg_ALUOP=0;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b001010:      //slti
            begin
                Reg_ALUOP=11;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b001011:      //sltiu
            begin
                Reg_ALUOP=4;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b001000:      //addi
            begin
                Reg_ALUOP=9;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b001001:      //addiu
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b001111:      //lui
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b000100:      // beq
            begin
                Reg_ALUOP=0;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b000101:      // bne
            begin
                Reg_ALUOP=0;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b000001:      //bgez & bltz
            begin
                Reg_ALUOP=0;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b000111:      //bgtz
            begin
                Reg_ALUOP=0;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b000110:      //blez
            begin
                Reg_ALUOP=0;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b100011:      //lw
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b100000:   //lb
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b100100:   //lbu
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b100001:   //lh
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b100101:   //lhu
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b101011:      //sw
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b101000:    //sb
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b101001:    //sh
            begin
                Reg_ALUOP=2;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        6'b000011:      //jal
            begin
                Reg_ALUOP=0;
                Reg_ALUSrc=1;
                RegDst=2;
            end
		  6'b000010:      //j
            begin
                Reg_ALUOP=0;
                Reg_ALUSrc=1;
                RegDst=0;       //change
            end
          6'b010000:      //mfc0
            begin
                if ({Instr_in[5:0]}==6'b011000) begin
                    Reg_ALUOP=0;
                    Reg_ALUSrc=1;
                    RegDst=0;
                end
                else begin
                    if({Instr_in[25:21]}==5'b00000) begin       //mfc0
                        Reg_ALUOP=0;
                        Reg_ALUSrc=1;
                        RegDst=0;
                    end
                    else begin                                  //mtc0
                        Reg_ALUOP=0;
                        Reg_ALUSrc=1;
                        RegDst=0;
                    end
                end
            end
        6'b000000:
            begin
                case (Instr_in[5:0])
                    6'b010000:       //mfhi
                        begin
                           Reg_ALUOP=0;
                           Reg_ALUSrc=1;
                           RegDst=1;
                        end
                    6'b010010:       //mflo
                        begin
                           Reg_ALUOP=0;
                           Reg_ALUSrc=1;
                           RegDst=1;
                        end
                    6'b010001:       //mthi
                        begin
                           Reg_ALUOP=0;
                           Reg_ALUSrc=1;
                           RegDst=0;
                        end
                    6'b010011:       //mtlo
                        begin
                           Reg_ALUOP=0;
                           Reg_ALUSrc=1;
                           RegDst=0;
                        end
                    6'b100001:      //addu
                        begin
                            Reg_ALUOP=2;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b100000:      //add
                        begin
                            Reg_ALUOP=9;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b000011:   //sra算术
                        begin
                            Reg_ALUOP=15;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b000010:   //srl逻辑
                        begin
                            Reg_ALUOP=14;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b000100:      //sllv
                        begin
                            Reg_ALUOP=7;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b000110:      //srlv
                        begin
                            Reg_ALUOP=5;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b000111:      //srav
                        begin
                            Reg_ALUOP=12;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b101010:     //slt
                        begin
                            Reg_ALUOP=11;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b101011:     //sltu
                        begin
                            Reg_ALUOP=4;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b100011:      //subu
                        begin
                            Reg_ALUOP=6;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b100010:      //sub
                        begin
                            Reg_ALUOP=10;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b100101:      //or
                        begin
                            Reg_ALUOP=1;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b100100:      //and
                        begin
                            Reg_ALUOP=0;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b100110:      //xor
                        begin
                            Reg_ALUOP=3;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b100111:      //nor
                        begin
                            Reg_ALUOP=8;
                            Reg_ALUSrc=0;
                            RegDst=1;
                        end
                    6'b001000:      //jr
                        begin
                            Reg_ALUOP=0;
                            Reg_ALUSrc=1;
                            RegDst=0;
                        end
                    6'b001001:     //jalr
                        begin
                            Reg_ALUOP=0;
                            Reg_ALUSrc=1;
                            RegDst=1;
                        end
                    6'b000000:      //nop & sll
                        begin
                            if(Instr_in==32'b0)  //nop
                            begin
                                Reg_ALUOP=0;
                                Reg_ALUSrc=1;
                                RegDst=0;
                            end
                            else begin          //sll
                                Reg_ALUOP=13;
                                Reg_ALUSrc=0;
                                RegDst=1;
                            end
                        end
                    6'b011000:       //mult
                        begin
                           Reg_ALUOP=0;
                           Reg_ALUSrc=1;
                           RegDst=0;
                        end
                    6'b011001:       //multu
                        begin
                           Reg_ALUOP=0;
                           Reg_ALUSrc=1;
                           RegDst=0;
                        end
                    6'b011010:       //div
                        begin
                           Reg_ALUOP=0;
                           Reg_ALUSrc=1;
                           RegDst=0;
                        end
                    6'b011011:       //divu
                        begin
                           Reg_ALUOP=0;
                           Reg_ALUSrc=1;
                           RegDst=0;
                        end
                    default:
                        begin
                            Reg_ALUOP=0;
                            Reg_ALUSrc=1;
                            RegDst=0;
                        end
                endcase
            end
            default:
            begin
                Reg_ALUOP=0;
                Reg_ALUSrc=1;
                RegDst=0;
            end
        endcase
    end

endmodule
